module select_freq (
  input reset,
  input 
);

endmodule